// =============================================================================
// audrey_top_test.sv
// Audrey — First Audio Test Top Level
//
// Project : rexta / Audrey
// Device  : Tang Nano 1K (Gowin GW1NZ-LV1)
// Author  : rexta project
// Version : 0.2
//
// Hardwired single voice driving PCM5102A via I2S.
// No SPI, no register file — just a fixed note to verify the audio chain.
//
// Hardwired voice settings:
//   Waveform  : Sawtooth
//   Frequency : ~440Hz (middle A)
//   ADSR      : fast attack, full sustain, gate always on
//
// Clock:
//   27MHz oscillator on pin 47.
//   Gowin rPLL generates 48.6MHz audio clock.
//   Sample rate: 48.6MHz / 32 / 32 = 47.46kHz (~1% flat, fine for testing)
//   Frequency word for 440Hz at 47.46kHz:
//     freq = round(440 * 65536 / 47460) = 0x0261
//
// PCM5102A breakout connections:
//   BCK  <- i2s_bclk  (pin 22)
//   DIN  <- i2s_data  (pin 23)
//   LCK  <- i2s_lrclk (pin 24)
//   SCK  <- leave floating (internal PLL)
//   XSMT <- VCC (unmute — must be high!)
//   GND  <- GND
//   VCC  <- 3.3V
// =============================================================================

module audrey_top_test (
    input  logic clk_27m,       // 27MHz oscillator (pin 47)

    // I2S output to PCM5102A
    output logic i2s_bclk,
    output logic i2s_lrclk,
    output logic i2s_data,

    // RGB LED (active low)
    output logic led_r,
    output logic led_g,
    output logic led_b,

    // Debug
    output logic dbg_req
);

// =============================================================================
// PLL — 27MHz -> 48.6MHz
// Generated by Gowin IP Core Generator (rPLL)
// =============================================================================
logic clk_audio;
logic pll_locked;

Gowin_rPLL pll (
    .clkin  (clk_27m),
    .clkout (clk_audio)
);

// lock port not enabled in PLL IP - tied high
// To add: regenerate Gowin_rPLL with lock output checked in IP Core Generator
assign pll_locked = 1'b1;

// =============================================================================
// Reset — hold for 256 cycles after PLL locks
// =============================================================================
logic [7:0] reset_counter;
logic       rst_n;

always @(posedge clk_audio) begin
    if (!pll_locked) begin
        reset_counter <= 8'h0;
        rst_n         <= 1'b0;
    end else if (!rst_n) begin
        if (reset_counter == 8'hFF)
            rst_n <= 1'b1;
        else
            reset_counter <= reset_counter + 8'h1;
    end
end

// =============================================================================
// I2S transmitter
// =============================================================================
logic        sample_req;
logic [15:0] left_sample;
logic [15:0] right_sample;

i2s_tx i2s (
    .clk        (clk_audio),
    .rst_n      (rst_n),
    .left_in    (left_sample),
    .right_in   (right_sample),
    .sample_req (sample_req),
    .bclk       (i2s_bclk),
    .lrclk      (i2s_lrclk),
    .data       (i2s_data)
);

// =============================================================================
// Voice engine — single hardwired voice
// Sawtooth, gate always on, ~440Hz
// =============================================================================
logic [15:0] voice_sample;

wavegen voice (
    .clk          (clk_audio),
    .rst_n        (rst_n),
    .sample_strobe(sample_req),

    .wave_ctrl    (8'b0000_1001),   // SAW=1, GATE=1
    .freq         (16'h0261),       // ~440Hz at 47.46kHz sample rate
    .pulse_width  (12'h800),        // 50% (unused for saw)

    .attack       (4'd1),           // 8ms attack
    .decay        (4'd0),           // minimal decay
    .sustain      (4'd15),          // full sustain
    .release_rate (4'd3),           // 72ms release

    .next_msb     (1'b0),
    .next_sync    (1'b0),
    .this_msb     (),
    .this_sync    (),

    .sample_out   (voice_sample)
);

// Mono — same sample to both channels
assign left_sample  = voice_sample;
assign right_sample = voice_sample;

// Debug output
assign dbg_req = sample_req;

// =============================================================================
// RGB LED — green heartbeat, others off
// Active low
// =============================================================================
logic [25:0] led_counter;
always @(posedge clk_audio) begin
    if (!rst_n)
        led_counter <= 26'h0;
    else
        led_counter <= led_counter + 26'h1;
end

assign led_r = 1'b1;                // off
assign led_g = ~led_counter[25];    // heartbeat ~0.7Hz
assign led_b = 1'b1;                // off

endmodule