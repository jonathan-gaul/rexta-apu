module apu_top (
);



endmodule